Current Feedback Amplifier

** Including necessary files **
.include OPAMP.MOD

** Defining parameters for output **
.CSPARAM RF=10k
.CSPARAM RL=10k

** Circuit Description **
I1 0 N1 1m
RF N1 N2 10k
RM N2 0 100
RL N2 N4 10k
XU2 0 N1 N4 OPAMP1

** Analysis Request **
.tran 0.1 10

** Output Request **
.control

run
* If = (V(N1) - V(N2))/RF
* Is = 1m
* Io = (V(N2) - V(N4))/RL

wrdata ep18btech11016_feed_gain.dat (V(N1) - V(N2))/(V(N2) - V(N4))
wrdata ep18btech11016_cl_gain.dat (V(N2) - V(N4))/(RL*1m)
.endc
.end
